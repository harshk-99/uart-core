`ifndef UART_ENV_PKG
`define UART_ENV_PKG

package uart_env_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

//////////////////////////////////////////////////////////
// importing packages : agent,ref model, register ...
/////////////////////////////////////////////////////////
  
import uart_agent_pkg::*;

//////////////////////////////////////////////////////////
// include top env files /////////////////////////////////
//////////////////////////////////////////////////////////

`include "uart_scoreboard.sv"
`include "uart_env.sv"

endpackage
`endif
